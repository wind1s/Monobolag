library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity uMem is
  port (
    Address : in unsigned(6 downto 0);
    Data : out std_logic_vector(25 downto 0)
  );
end entity;

architecture Behavioral of uMem is

-- micro Memory
type u_mem_t is array (0 to 127) of std_logic_vector(25 downto 0);
constant u_mem_c : u_mem_t :=
   --      OP TDB FDB TAB  P LC  SEQ    uADR 
  (
  0 =>  b"0000_000_000_011_01_0000_0000000",  -- Hämtfas
  1 =>  b"0000_000_000_000_00_0011_0000000",
  2 =>  b"0000_001_101_000_00_0010_0000000",  -- Omedelbar; K2 prolog
  3 =>  b"0000_110_101_000_00_0010_0000000",  -- Direkt register; K2 prolog
  4 =>  b"0000_010_101_001_00_0010_0000000",  -- Direkt till/från; K2 prolog
  5 =>  b"0000_010_101_110_00_0010_0000000",  -- Indirekt till/från; K2 prolog
  6 =>  b"0010_000_000_000_00_0000_0000000",  -- Indexerad till/från; K2 prolog
  7 =>  b"0000_010_101_100_00_0010_0000000",
  8 =>  b"0000_101_110_000_00_0001_0000000",  -- Omedelbar, Direkt register, Direkt/indirekt/indexerad från; K3
  9 =>  b"0000_101_010_001_00_0001_0000000",  -- Direkt till; K3
  10 => b"0000_101_010_110_00_0001_0000000", -- Indirekt till; K3
  11 => b"0010_000_000_000_00_0000_0000000", -- Indexerad till; K3
  12 => b"0000_101_010_100_00_0001_0000000",
  13 => b"0000_000_000_000_00_0001_0000000", -- NOP
  14 => b"0000_000_000_000_00_1111_0000000", -- HALT
  15 => b"0000_101_011_000_00_0001_0000000", -- JMP
  16 => b"1101_101_000_000_00_0000_0000000", -- MOV
  17 => b"0000_100_101_000_00_0100_0000000", -- SAVE AR
  18 => b"0011_101_000_000_00_0101_0010001", -- ADD
  19 => b"0100_101_000_000_00_0101_0010001", -- SUB
  20 => b"0101_101_000_000_00_0101_0010001", -- MUL
  21 => b"1011_101_000_000_00_0101_0010001", -- INC
  22 => b"1100_101_000_000_00_0101_0010001", -- DEC
  23 => b"0110_101_000_000_00_0101_0010001", -- AND
  24 => b"0111_101_000_000_00_0101_0010001", -- OR
  25 => b"1000_101_000_000_00_0101_0010001", -- XOR
  26 => b"0100_101_000_000_00_0001_0000000", -- CMP
  27 => b"0001_000_000_000_00_0101_0010001", -- CLR
  28 => b"0000_011_010_010_11_0000_0000000", -- CALL
  29 => b"0000_101_011_000_00_0001_0000000",
  30 => b"0000_000_000_000_10_0000_0000000", -- RET
  31 => b"0000_010_011_010_00_0001_0000000",
  32 => b"0000_101_010_010_11_0001_0000000", -- PUSH
  33 => b"0000_000_000_000_10_0000_0000000", -- POP
  34 => b"0000_010_101_010_00_0100_0000000", 
  35 => b"0000_000_000_000_00_0111_0001111", -- JEQ
  36 => b"0000_000_000_000_00_0001_0000000",
  37 => b"0000_000_000_000_00_0110_0001111", -- JNE
  38 => b"0000_000_000_000_00_0001_0000000",
  39 => b"0000_000_000_000_00_0111_0000000", -- JGT
  40 => b"0000_000_000_000_00_1100_0101011", -- JGE
  41 => b"0000_000_000_000_00_1010_0001111", -- LABEL V0
  42 => b"0000_000_000_000_00_0001_0000000",
  43 => b"0000_000_000_000_00_1011_0001111", -- LABEL v1
  44 => b"0000_000_000_000_00_0001_0000000",
  45 => b"0000_000_000_000_00_0111_0001111", -- JLE
  46 => b"0000_000_000_000_00_1100_0101001", -- JLT
  47 => b"0000_000_000_000_00_0101_0101011",
  48 => b"0000_000_000_000_00_1001_0001111", -- JCS
  49 => b"0000_000_000_000_00_0001_0000000",
  50 => b"1001_101_000_000_00_0101_0010001", -- LSL
  51 => b"1010_101_000_000_00_0101_0010001", -- LSR
  52 => b"0000_000_000_000_00_0110_0000000", -- MOVZ
  53 => b"0000_000_000_000_00_0101_0010000",
  54 => b"0000_000_000_000_00_0110_0000000", -- ADDZ
  55 => b"0000_000_000_000_00_0101_0010010", 
  56 => b"0000_000_000_000_00_0110_0000000", -- MULZ
  57 => b"0000_000_000_000_00_0101_0010100",
  58 => b"0000_000_000_000_00_0110_0000000", -- ANDZ
  59 => b"0000_000_000_000_00_0101_0010111",
  60 => b"0000_000_000_000_00_0110_0000000", -- ORZ
  61 => b"0000_000_000_000_00_0101_0011000",
  others => b"0000_000_000_000_00_1111_0000000" -- HALT om vi hamnar på konstig address.
  );

signal u_mem : u_mem_t := u_mem_c;

begin
  Data <= u_mem(to_integer(Address));

end Behavioral;
